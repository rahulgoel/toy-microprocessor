----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:23:35 03/31/2012 
-- Design Name: 
-- Module Name:    aftrinp - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity aftrinp1 is
    Port ( bitmodeout44 : in  STD_LOGIC_VECTOR (3 downto 0);
           bitreg1out22 : in  STD_LOGIC_VECTOR (1 downto 0);
           bitreg2out22 : in  STD_LOGIC_VECTOR (1 downto 0);
			  bitintout88: in STD_LOGIC_VECTOR (7 downto 0);
			  --out_port1 : out STD_LOGIC_VECTOR (7 downto 0);
			  clk :in std_logic;
			 --out_port2: out STD_LOGIC;
			 stack_out :out STD_LOGIC_VECTOR (7 downto 0);
			  oreg0,oreg1,oreg2,oreg3 : out STD_LOGIC_VECTOR (7 downto 0);
			 jumpp1: out STD_LOGIC_VECTOR (7 downto 0) );
			  
end aftrinp1;


architecture Behavioral of aftrinp1 is

signal treg1,treg2,reg0,reg1,reg2,reg3,temp1,Data_out,stack_ptr1,jmp_stk,jmp_stk_t : STD_LOGIC_VECTOR (7 downto 0);
shared variable var88: Std_logic_vector(7 downto 0);

				
--variable shift:STD_LOGIC:='0';
signal PUSH_barPOP , shift:STD_LOGIC;
--type mem_type is array (255 downto 0) of std_logic_vector(7 downto 0);
--signal stack_mem : mem_type := (others => (others => '0'));
shared variable stack_ptr : integer := 255;
signal full,empty : std_logic := '0'; 

function memory(add : std_logic_vector(7 downto 0)) return std_logic_vector is
variable ret :std_logic_vector(7 downto 0);
variable index :integer;
type dataout is array (0 to 255) of STD_LOGIC_VECTOR (7 downto 0);
variable arr: dataout;

begin

arr(0):=('0','0','1','0','0','0','0','1');
arr(1):=('1','1','0','1','1','0','1','0');
arr(2):=('1','0','1','1','0','1','0','1');
arr(3):=('1','1','0','0','0','1','0','1');
arr(4):=('0','1','0','1','1','0','0','1');
arr(5):=('1','0','1','0','0','1','0','1');
arr(6):=('0','1','0','0','1','1','0','1');
arr(7):=('0','0','1','1','1','1','0','1');
arr(8):=('1','0','1','1','0','1','0','1');
arr(9):=('1','0','1','0','0','0','1','1');
arr(10):=('1','0','1','0','0','1','1','1');
arr(11):=('1','0','1','1','0','0','0','1');
arr(12):=('0','0','1','1','1','0','1','1');
arr(13):=('1','0','1','0','0','0','1','1');
arr(14):=('1','0','1','0','1','0','1','1');
arr(15):=('0','1','1','0','1','0','1','1');
arr(16):=('0','1','1','0','0','0','0','1');
arr(17):=('0','1','1','0','1','1','0','1');
arr(18):=('1','0','1','1','0','1','0','1');
arr(19):=('0','0','1','1','0','1','0','1');
arr(20):=('0','1','1','0','0','1','0','0');
arr(21):=('1','1','1','1','1','0','0','0');
arr(22):=('1','1','1','0','0','0','0','0');
arr(23):=('0','1','1','1','0','0','1','1');
arr(24):=('0','0','1','0','0','0','1','1');
arr(25):=('0','0','1','1','0','0','1','1');
arr(26):=('0','0','1','1','0','1','0','1');
arr(27):=('1','0','1','0','0','1','0','1');
arr(28):=('1','0','1','0','0','0','1','1');
arr(29):=('0','0','1','1','0','0','1','1');
arr(30):=('0','0','1','1','1','0','0','1');
arr(31):=('0','1','1','0','1','0','0','1');
arr(32):=('0','1','1','0','1','0','0','0');
arr(33):=('0','0','1','0','0','1','0','0');
arr(34):=('0','1','0','0','0','1','0','1');
arr(35):=('0','0','0','0','1','0','0','1');
arr(36):=('0','0','1','0','1','1','1','1');
arr(37):=('1','0','1','0','1','0','1','1');
arr(38):=('1','1','1','0','0','0','0','1');
arr(39):=('0','1','1','0','1','0','0','1');
arr(40):=('0','0','1','0','1','1','0','1');
arr(41):=('0','0','1','0','0','1','1','1');
arr(42):=('0','0','1','0','1','0','1','1');
arr(43):=('0','0','1','0','1','0','0','1');
arr(44):=('1','0','1','0','1','0','0','1');
arr(45):=('1','1','1','0','0','0','0','1');
arr(46):=('0','1','1','0','1','0','0','1');
arr(47):=('0','0','1','0','1','0','1','1');
arr(48):=('0','0','1','0','0','0','1','1');
arr(49):=('0','1','1','0','0','0','1','0');
arr(50):=('0','1','1','1','0','0','0','1');
arr(51):=('0','0','1','1','1','0','0','1');
arr(52):=('0','1','1','0','1','0','0','1');
arr(53):=('0','0','0','1','0','0','1','1');
arr(54):=('1','0','1','0','0','1','1','1');
arr(55):=('1','1','1','0','1','0','0','1');
arr(56):=('0','0','1','0','1','0','0','1');
arr(57):=('0','1','0','0','0','0','0','1');
arr(58):=('0','1','1','1','1','0','0','0');
arr(59):=('0','0','1','1','0','0','1','0');
arr(60):=('0','0','0','1','1','0','0','1');
arr(61):=('1','0','0','0','0','0','0','1');
arr(62):=('1','0','1','0','0','1','0','1');
arr(63):=('0','0','1','0','0','1','1','1');
arr(64):=('1','0','1','0','0','0','0','0');
arr(65):=('1','0','1','0','0','0','0','1');
arr(66):=('0','1','1','0','0','0','0','1');
arr(67):=('0','0','1','1','0','1','0','1');
arr(68):=('0','0','1','1','0','1','0','1');
arr(69):=('0','0','1','0','0','0','1','1');
arr(70):=('1','0','1','0','0','1','1','1');
arr(71):=('0','1','0','0','0','1','0','1');
arr(72):=('0','1','1','0','0','1','0','1');
arr(73):=('0','0','0','0','1','0','0','1');
arr(74):=('1','0','1','0','0','0','1','0');
arr(75):=('1','0','1','1','0','1','0','1');
arr(76):=('0','0','1','1','0','1','0','1');
arr(77):=('1','1','1','0','0','0','0','1');
arr(78):=('0','0','1','0','0','1','1','0');
arr(79):=('1','1','1','0','1','1','0','1');
arr(80):=('0','1','1','0','0','1','0','1');
arr(81):=('0','0','1','0','0','1','1','1');
arr(82):=('1','0','1','0','0','0','1','0');
arr(83):=('0','1','1','0','0','0','0','1');
arr(84):=('0','0','1','1','1','0','1','1');
arr(85):=('0','0','1','0','0','0','0','1');
arr(86):=('0','0','1','0','1','0','1','1');
arr(87):=('0','0','1','0','1','0','0','1');
arr(88):=('1','1','1','0','1','0','0','1');
arr(89):=('0','1','1','0','1','0','0','1');
arr(90):=('0','0','1','0','1','0','0','1');
arr(91):=('0','0','1','1','0','0','0','1');
arr(92):=('1','0','0','1','0','0','0','1');
arr(93):=('1','0','0','0','0','1','0','1');
arr(94):=('0','0','0','0','0','0','0','1');
arr(95):=('1','1','1','0','0','0','0','1');
arr(96):=('0','1','1','1','0','1','0','1');
arr(97):=('1','0','1','0','1','1','0','1');
arr(98):=('1','0','1','0','0','1','0','1');
arr(99):=('0','0','1','0','1','1','0','0');
arr(100):=('1','0','1','0','0','1','0','1');
arr(101):=('1','1','1','0','1','0','0','1');
arr(102):=('0','0','1','0','1','0','1','1');
arr(103):=('0','1','1','0','0','1','0','1');
arr(104):=('0','1','1','0','0','1','0','1');
arr(105):=('1','1','1','0','0','0','0','0');
arr(106):=('0','1','1','1','0','0','1','1');
arr(107):=('1','1','1','0','0','0','1','1');
arr(108):=('0','1','0','0','0','0','0','1');
arr(109):=('1','0','0','0','0','1','1','1');
arr(110):=('0','0','1','1','0','1','0','1');
arr(111):=('0','1','1','0','0','0','1','0');
arr(112):=('0','1','0','0','0','0','1','1');
arr(113):=('1','0','0','0','0','1','1','1');
arr(114):=('1','0','1','1','0','0','1','0');
arr(115):=('1','0','1','0','1','0','0','1');
arr(116):=('1','0','0','0','1','0','0','1');
arr(117):=('0','1','1','0','1','1','1','1');
arr(118):=('0','1','1','0','1','0','0','1');
arr(119):=('1','0','0','0','1','0','0','1');
arr(120):=('1','1','0','0','0','0','1','1');
arr(121):=('0','0','1','0','1','0','1','1');
arr(122):=('1','0','0','1','0','0','0','1');
arr(123):=('0','1','1','0','1','1','0','1');
arr(124):=('1','0','1','0','0','1','0','1');
arr(125):=('1','0','1','0','1','1','0','0');
arr(126):=('0','1','1','0','0','0','0','0');
arr(127):=('0','1','1','0','0','0','1','1');
arr(128):=('1','0','1','0','1','0','0','1');
arr(129):=('1','0','1','0','1','0','0','0');
arr(130):=('0','0','1','1','0','0','1','0');
arr(131):=('0','0','1','1','0','1','1','1');
arr(132):=('0','0','1','0','0','1','1','1');
arr(133):=('0','1','1','0','1','0','0','1');
arr(134):=('0','1','1','1','0','0','0','1');
arr(135):=('0','0','1','1','0','0','0','0');
arr(136):=('0','1','1','1','0','0','0','1');
arr(137):=('0','1','1','0','0','0','1','1');
arr(138):=('0','0','1','0','1','0','1','1');
arr(139):=('0','0','1','0','0','1','0','1');
arr(140):=('0','0','1','0','0','1','0','1');
arr(141):=('1','0','1','1','0','0','0','0');
arr(142):=('1','1','0','1','0','0','0','1');
arr(143):=('0','0','1','0','1','0','0','0');
arr(144):=('1','1','0','0','1','0','0','1');
arr(145):=('0','1','0','0','0','0','1','0');
arr(146):=('0','0','0','0','1','1','1','1');
arr(147):=('0','0','0','0','0','1','1','1');
arr(148):=('1','1','1','0','0','1','1','1');
arr(149):=('0','0','1','1','0','1','0','0');
arr(150):=('0','0','1','0','1','1','0','1');
arr(151):=('1','1','1','0','1','0','0','1');
arr(152):=('0','1','1','0','1','0','0','1');
arr(153):=('0','0','1','0','1','0','0','1');
arr(154):=('0','0','0','0','1','1','0','1');
arr(155):=('0','0','1','1','0','0','0','1');
arr(156):=('0','0','1','1','0','0','1','0');
arr(157):=('0','0','1','0','0','0','1','1');
arr(158):=('1','0','1','0','0','0','1','1');
arr(159):=('0','1','1','0','0','0','0','1');
arr(160):=('0','1','1','0','0','0','0','1');
arr(161):=('0','0','0','0','0','0','0','1');
arr(162):=('0','0','1','1','0','0','0','1');
arr(163):=('0','0','1','1','1','0','0','1');
arr(164):=('0','0','1','0','1','0','0','1');
arr(165):=('0','0','1','1','1','0','0','0');
arr(166):=('0','0','0','0','1','0','0','1');
arr(167):=('0','0','1','0','1','0','0','0');
arr(168):=('0','0','1','0','0','0','1','0');
arr(169):=('1','0','1','0','0','0','1','1');
arr(170):=('1','0','1','0','0','0','0','1');
arr(171):=('1','1','1','0','0','0','0','1');
arr(172):=('0','0','1','1','0','0','0','1');
arr(173):=('0','0','1','0','1','0','0','1');
arr(174):=('0','0','1','0','0','1','0','1');
arr(175):=('0','0','1','0','0','1','1','0');
arr(176):=('0','0','1','0','0','0','0','1');
arr(177):=('1','0','1','0','0','0','0','0');
arr(178):=('1','0','1','0','0','0','0','1');
arr(179):=('1','0','1','1','0','1','0','1');
arr(180):=('0','0','1','1','1','0','0','1');
arr(181):=('0','0','1','0','1','1','0','1');
arr(182):=('0','0','1','1','0','1','0','1');
arr(183):=('0','0','1','1','1','0','0','1');
arr(184):=('1','0','1','0','1','0','0','1');
arr(185):=('1','1','0','0','0','0','0','1');
arr(186):=('0','0','0','0','1','0','0','0');
arr(187):=('0','0','1','0','0','1','1','1');
arr(188):=('0','0','1','1','0','1','0','1');
arr(189):=('0','0','1','1','0','0','0','1');
arr(190):=('0','0','1','0','0','0','0','1');
arr(191):=('0','0','1','1','0','1','0','1');
arr(192):=('0','1','1','0','0','1','0','1');
arr(193):=('0','1','0','0','0','0','0','0');
arr(194):=('0','0','1','0','1','1','0','0');
arr(195):=('0','0','1','0','1','1','0','1');
arr(196):=('0','0','1','0','0','1','0','0');
arr(197):=('0','0','1','0','0','1','0','0');
arr(198):=('0','0','1','1','0','1','1','1');
arr(199):=('0','0','1','0','1','0','0','1');
arr(200):=('0','1','1','0','0','1','0','1');
arr(201):=('0','1','1','0','0','0','0','1');
arr(202):=('1','1','1','0','0','0','0','1');
arr(203):=('1','0','1','0','1','0','0','1');
arr(204):=('0','0','1','1','1','0','0','1');
arr(205):=('0','1','0','0','0','0','0','1');
arr(206):=('1','0','1','0','0','0','0','1');
arr(207):=('0','0','1','0','0','0','0','1');
arr(208):=('0','1','1','0','0','0','0','1');
arr(209):=('0','0','1','1','0','0','0','1');
arr(210):=('0','0','1','0','1','0','0','1');
arr(211):=('0','0','1','0','0','1','0','1');
arr(212):=('0','0','1','0','0','0','0','1');
arr(213):=('0','0','1','0','0','0','1','1');
arr(214):=('0','0','1','1','0','0','1','1');
arr(215):=('0','0','1','0','0','0','0','1');
arr(216):=('0','0','1','0','1','1','1','1');
arr(217):=('0','0','1','0','1','0','0','1');
arr(218):=('0','0','1','0','1','0','0','1');
arr(219):=('0','0','1','1','0','0','0','1');
arr(220):=('0','0','0','0','0','0','0','0');
arr(221):=('0','0','1','0','0','1','0','0');
arr(222):=('0','0','1','0','1','1','0','1');
arr(223):=('0','1','1','0','1','0','0','1');
arr(224):=('0','1','0','1','0','0','0','1');
arr(225):=('0','0','1','0','1','1','0','1');
arr(226):=('0','0','0','0','1','0','1','1');
arr(227):=('0','0','0','0','0','0','0','1');
arr(228):=('0','1','0','0','0','0','0','1');
arr(229):=('1','0','1','0','0','0','0','1');
arr(230):=('1','1','1','0','0','0','0','1');
arr(231):=('0','1','1','0','0','0','0','1');
arr(232):=('0','1','1','1','0','0','0','1');
arr(233):=('0','0','1','0','0','1','0','1');
arr(234):=('0','0','1','0','1','0','0','1');
arr(235):=('0','0','1','0','0','1','0','1');
arr(236):=('0','0','1','0','0','1','1','0');
arr(237):=('0','0','1','0','0','0','0','0');
arr(238):=('0','0','1','0','0','0','1','0');
arr(239):=('0','0','0','0','0','0','1','1');
arr(240):=('0','0','0','0','0','0','0','1');
arr(241):=('0','0','1','1','0','0','0','1');
arr(242):=('0','0','0','0','0','0','0','1');
arr(243):=('0','0','1','1','0','0','0','1');
arr(244):=('0','0','1','0','0','1','1','1');
arr(245):=('0','0','1','0','0','1','0','1');
arr(246):=('0','0','1','0','0','0','1','1');
arr(247):=('0','0','1','1','0','0','0','1');
arr(248):=('0','0','1','0','0','0','0','1');
arr(249):=('0','0','0','0','0','0','0','1');
arr(250):=('0','0','1','1','0','0','0','1');
arr(251):=('0','1','0','0','0','0','0','1');
arr(252):=('0','0','1','0','0','0','0','1');
arr(253):=('0','0','1','0','0','0','0','1');
arr(254):=('1','1','1','0','0','0','0','1');
arr(255):=('1','0','1','0','0','0','0','1');

index := conv_integer(unsigned(add));

ret:=arr(index);
return ret;
end;


type stack is array (255 downto 0) of std_logic_vector(7 downto 0);
--signal stack_mem : mem_type := (others => (others => '0'));

 function stock(temp1: std_logic_vector(7 downto 0);
					shift: std_logic
					) return std_logic_vector is
variable stock_out : std_logic_vector(7 downto 0);
variable stack1:stack;
--variable s : line ;
begin
	
	--if (rising_edge(clk)) then
	
		if shift = '1' and stack_ptr /= 0 then
		stack1(stack_ptr) := temp1;
		stack_ptr := stack_ptr -1 ;
		stock_out := temp1;
		end if;
		
		if shift = '0' and stack_ptr /= 255 then
		stock_out := stack1(stack_ptr);
		stack_ptr := stack_ptr + 1 ;
		elsif shift = '0' and stack_ptr = 255 then
		--write(s, "Stack is empty");
		end if;
		
	--end if;
	return stock_out;
end function stock;

begin
--procedure stack( signal temp1 : in std_logic_vector (7 downto 0);
	--				  signal shift : in std_logic;
		--				signal clk	: in std_logic );
--		begin
--		
--		if (rising edge(clk)) then
		
--		if shift = '1' and full = '0' then
			--stack_mem(stack_ptr) <= temp1;
			--stack_out<=stack_mem(stack_ptr);	
		
--			if(stack_ptr /= 0) then
 --               stack_ptr <= stack_ptr - 1;
--         end if;
			 --setting full and empty flags
--         if(stack_ptr = 0) then
--                full <= '1';
--                empty <= '0';
--         elsif(stack_ptr = 255) then
--                full <= '0';
--                empty <= '1';
--         else
--                full <= '0';
--                empty <= '0';
--         end if;
--		end if;
		
--		if shift = '0' and empty = '0' then
--			if(stack_ptr /= 255) then   
--                Data_Out <= stack_mem(stack_ptr); 
--                stack_ptr <= stack_ptr + 1;
--			end if ; 
            --setting full and empty flags
--         if(stack_ptr = 0) then
--                full <= '1';
--                empty <= '0';
--         elsif(stack_ptr = 255) then
--                full <= '0';
--                empty <= '1';
--         else
--                full <= '0';
--                empty <= '0';
--			end if;
--		end if;
		
--		end if
		
--		end procedure stack ;

reg0<="10100010";--162
reg1<="11111010";--250
reg2<="10111010";--192
reg3<="10101010";--180



process(bitmodeout44, bitreg1out22, bitreg2out22, bitintout88,clk)


begin
oreg0<="10100010";--162
oreg1<="11111010";--250
oreg2<="10111010";--192
oreg3<="10101010";--180
jmp_stk<="00000000";
--bitreg2out2 <= "00" ;
--register 1 value

case bitreg1out22 is
when "00"=>treg1<=reg0;
when "01"=>treg1<=reg1;
when "10"=>treg1<=reg2;
when "11"=>treg1<=reg3;
when others => reg3 <= treg1;
end case;
-- register 2 value
case bitreg2out22 is
when "00"=>treg2<=reg0;
when "01"=>treg2<=reg1;
when "10"=>treg2<=reg2;
when "11"=>treg2<=reg3;
when others => reg3 <= treg1;
end case;


--modes statement
if(bitmodeout44="0000") then
treg1<=treg2;

case bitreg1out22 is
when "00"=>oreg0<=treg1;
when "01"=>oreg1<=treg1;
when "10"=>oreg2<=treg1;
when "11"=>oreg3<=treg1;
when others => reg3 <= treg1;
end case;


elsif (bitmodeout44="0001")then
 treg1<=bitintout88;
 case bitreg1out22 is
when "00"=>oreg0<=treg1;
when "01"=>oreg1<=treg1;
when "10"=>oreg2<=treg1;
when "11"=>oreg3<=treg1;
when others => reg3 <= treg1;
end case;



elsif (bitmodeout44="0010")then
treg1<=treg1+treg2;
case bitreg1out22 is
when "00"=>oreg0<=treg1;
when "01"=>oreg1<=treg1;
when "10"=>oreg2<=treg1;
when "11"=>oreg3<=treg1;
when others => reg3 <= treg1;
end case;


elsif (bitmodeout44="0011")then
treg1<=treg1+ bitintout88 ;
case bitreg1out22 is
when "00"=>oreg0<=treg1;
when "01"=>oreg1<=treg1;
when "10"=>oreg2<=treg1;
when "11"=>oreg3<=treg1;
when others => reg3 <= treg1;
end case;

elsif (bitmodeout44="0100")then
treg1<=treg1-treg2;
case bitreg1out22 is
when "00"=>oreg0<=treg1;
when "01"=>oreg1<=treg1;
when "10"=>oreg2<=treg1;
when "11"=>oreg3<=treg1;
when others => reg3 <= treg1;
end case;

elsif (bitmodeout44="0101")then
treg1<=treg1-bitintout88;
case bitreg1out22 is
when "00"=>oreg0<=treg1;
when "01"=>oreg1<=treg1;
when "10"=>oreg2<=treg1;
when "11"=>oreg3<=treg1;
when others => reg3 <= treg1;
end case;
--
--elsif (bitmodeout44="1001")then
--
--		jmp_stk_t <=bitintout88;
--		jmp_stk <=jmp_stk_t;
--		stack_out<=stock(jmp_stk,'1');

--elsif (bitmodeout44="0111")then
--procedure stack(bitintout88, '1', clk);
--jmp_stk_t <=bitintout88;
--var88:=stock(jmp_stk,'0');
--stack_out<=var88;
--jmp_stk <=var88;

		

elsif(bitmodeout44="1000") then
--procedure stack ( bitintout8, '0', clk);		  
stack_out <= memory(bitintout88);

elsif (bitmodeout44="0110")then
jmp_stk_t <=bitintout88;
jmp_stk <=bitintout88;
stack_out<=stock(jmp_stk,'1');



elsif (bitmodeout44="1010")then

elsif (bitmodeout44="1011")then

elsif (bitmodeout44="1100")then

elsif (bitmodeout44="1101")then

elsif (bitmodeout44="1110")then

elsif (bitmodeout44="1111")then

end if;
jumpp1<=jmp_stk;
end process ;

end Behavioral;



